../../normal/src/top.sv