../../normal/src/noc.sv