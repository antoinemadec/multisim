../../normal/src/cpu.sv